/*
 *  PicoSoC - A simple example SoC using PicoRV32
 *
 *  Copyright (C) 2017  Clifford Wolf <clifford@clifford.at>
 *
 *  Permission to use, copy, modify, and/or distribute this software for any
 *  purpose with or without fee is hereby granted, provided that the above
 *  copyright notice and this permission notice appear in all copies.
 *
 *  THE SOFTWARE IS PROVIDED "AS IS" AND THE AUTHOR DISCLAIMS ALL WARRANTIES
 *  WITH REGARD TO THIS SOFTWARE INCLUDING ALL IMPLIED WARRANTIES OF
 *  MERCHANTABILITY AND FITNESS. IN NO EVENT SHALL THE AUTHOR BE LIABLE FOR
 *  ANY SPECIAL, DIRECT, INDIRECT, OR CONSEQUENTIAL DAMAGES OR ANY DAMAGES
 *  WHATSOEVER RESULTING FROM LOSS OF USE, DATA OR PROFITS, WHETHER IN AN
 *  ACTION OF CONTRACT, NEGLIGENCE OR OTHER TORTIOUS ACTION, ARISING OUT OF
 *  OR IN CONNECTION WITH THE USE OR PERFORMANCE OF THIS SOFTWARE.
 *
 */

module hardware (
    input clk_16mhz,
    input pin_go,

    // onboard USB interface
    output pin_pu,
    output pin_usbp,
    output pin_usbn,

    // hardware UART
    output uart_out,
    input uart_in,

    output pin_7,
    output pin_8,


    // onboard SPI flash interface
    output flash_csb,
    output flash_clk,
    inout  flash_io0,
    inout  flash_io1,
    inout  flash_io2,
    inout  flash_io3
);
    assign pin_pu = 1'b1;
    assign pin_usbp = 1'b0;
    assign pin_usbn = 1'b0;

    wire clk = clk_16mhz;

    assign pin_8=clock_out[0];
  

    ///////////////////////////////////
    // Power-on Reset
    ///////////////////////////////////
    reg [5:0] reset_cnt = 0;
    wire resetn = &reset_cnt;

    always @(posedge clk) begin
        reset_cnt <= reset_cnt + !resetn;
    end

  
    ///////////////////////////////////
    // SPI Flash Interface
    ///////////////////////////////////
    wire flash_io0_oe, flash_io0_do, flash_io0_di;
    wire flash_io1_oe, flash_io1_do, flash_io1_di;
    wire flash_io2_oe, flash_io2_do, flash_io2_di;
    wire flash_io3_oe, flash_io3_do, flash_io3_di;

    SB_IO #(
        .PIN_TYPE(6'b 1010_01),
        .PULLUP(1'b 0)
    ) flash_io_buf [3:0] (
        .PACKAGE_PIN({flash_io3, flash_io2, flash_io1, flash_io0}),
        .OUTPUT_ENABLE({flash_io3_oe, flash_io2_oe, flash_io1_oe, flash_io0_oe}),
        .D_OUT_0({flash_io3_do, flash_io2_do, flash_io1_do, flash_io0_do}),
        .D_IN_0({flash_io3_di, flash_io2_di, flash_io1_di, flash_io0_di})
    );

    
  
    ///////////////////////////////////
    // Peripheral Bus
    ///////////////////////////////////
    wire        iomem_valid;
    reg         iomem_ready;
    wire [3:0]  iomem_wstrb;
    wire [31:0] iomem_addr;
    wire [31:0] iomem_wdata;
    reg [31:0] clock_out;
    reg  [31:0] iomem_rdata;

    reg [31:0] clockO=0;
    reg [31:0] gpio;
    reg [31:0] leds;

    reg writeEncoderL=0;
    reg writeEncoderR=0;
    wire [31:0] encoderValueL;
    wire [31:0] encoderValueR;
    reg [31:0] encoderDataL=0;
    reg [31:0] encoderDataR=0;
    

    reg[31:0] pinTest=0;
    assign pin_7=pinTest[0];

    always @(posedge clk) begin
        if (!resetn) begin
            gpio <= 0;
        end else begin
            iomem_ready <= 0;
            writeEncoderL <=0; 
            writeEncoderR <=0; 

            ///////////////////////////
            // GPIO Peripheral
            ///////////////////////////
            if (iomem_valid && !iomem_ready && iomem_addr[31:8] == 24'h030000) begin
                iomem_ready <= 1;
                iomem_rdata <= gpio;
                if (iomem_wstrb[0]) gpio[ 7: 0] <= iomem_wdata[ 7: 0];
                if (iomem_wstrb[1]) gpio[15: 8] <= iomem_wdata[15: 8];
                if (iomem_wstrb[2]) gpio[23:16] <= iomem_wdata[23:16];
                if (iomem_wstrb[3]) gpio[31:24] <= iomem_wdata[31:24];
            end

            if (iomem_valid && !iomem_ready && iomem_addr[31:8] == 24'h030001) begin
                iomem_ready <= 1;
                iomem_rdata <= pin_go;
                if (iomem_wstrb[0]) leds[ 7: 0] <= iomem_wdata[ 7: 0];
                if (iomem_wstrb[1]) leds[15: 8] <= iomem_wdata[15: 8];
                if (iomem_wstrb[2]) leds[23:16] <= iomem_wdata[23:16];
                if (iomem_wstrb[3]) leds[31:24] <= iomem_wdata[31:24];
                //leds=32'hffffffff;
            end

            if (iomem_valid && !iomem_ready && iomem_addr[31:8] == 24'h030002) begin
                iomem_ready <= 1;
                iomem_rdata <= clock_out;
                if (iomem_wstrb[0]) clockO[ 7: 0] <= iomem_wdata[ 7: 0];
                if (iomem_wstrb[1]) clockO[15: 8] <= iomem_wdata[15: 8];
                if (iomem_wstrb[2]) clockO[23:16] <= iomem_wdata[23:16];
                if (iomem_wstrb[3]) clockO[31:24] <= iomem_wdata[31:24];
            end

            if (iomem_valid && !iomem_ready && iomem_addr[31:8] == 24'h030009) begin
                iomem_ready <= 1;
                if (iomem_wstrb[0]) pinTest[ 7: 0] <= iomem_wdata[ 7: 0];
                if (iomem_wstrb[1]) pinTest[15: 8] <= iomem_wdata[15: 8];
                if (iomem_wstrb[2]) pinTest[23:16] <= iomem_wdata[23:16];
                if (iomem_wstrb[3]) pinTest[31:24] <= iomem_wdata[31:24];
            end
            
            ///////////////////////////
            // Template Peripheral
            ///////////////////////////
            if (iomem_valid && !iomem_ready && iomem_addr[31:24] == 8'h04) begin
                iomem_ready <= 1;
                iomem_rdata <= 32'h0;
            end
        end
    end

    ///////////////////////////////////
    // Custom Modules
    ///////////////////////////////////

    clock clock (
		.clk         (clk         ),
		.resetn      (resetn      ),
		.clock_out   (clock_out)
	);


    ///////////////////////////////////
    // PicoSOC
    ///////////////////////////////////

    picosoc #(
        .PROGADDR_RESET(32'h0005_0000), // beginning of user space in SPI flash
        .PROGADDR_IRQ(32'h0005_0010),
        .MEM_WORDS(2048)                // use 2KBytes of block RAM by default
    ) soc (
        .clk          (clk         ),
        .resetn       (resetn      ),

        .ser_tx       (uart_out       ),
        .ser_rx       (uart_in       ),

        .flash_csb    (flash_csb   ),
        .flash_clk    (flash_clk   ),

        .flash_io0_oe (flash_io0_oe),
        .flash_io1_oe (flash_io1_oe),
        .flash_io2_oe (flash_io2_oe),
        .flash_io3_oe (flash_io3_oe),

        .flash_io0_do (flash_io0_do),
        .flash_io1_do (flash_io1_do),
        .flash_io2_do (flash_io2_do),
        .flash_io3_do (flash_io3_do),

        .flash_io0_di (flash_io0_di),
        .flash_io1_di (flash_io1_di),
        .flash_io2_di (flash_io2_di),
        .flash_io3_di (flash_io3_di),

        .irq_5        (1'b0        ),
        .irq_6        (1'b0        ),
        .irq_7        (1'b0        ),

        .iomem_valid  (iomem_valid ),
        .iomem_ready  (iomem_ready ),
        .iomem_wstrb  (iomem_wstrb ),
        .iomem_addr   (iomem_addr  ),
        .iomem_wdata  (iomem_wdata ),
        .iomem_rdata  (iomem_rdata )
    );
endmodule