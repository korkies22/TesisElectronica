/*
 * Clock Module
 */

module pwm #(
	parameter DURATION_CYCLE=32
)(
	input clk,
    input resetn,
	input pwm_in,
	output pwm_out,
);
	reg [31:0] counterI=0;

    reg pwm_counter=0;

	reg [8:0] count_temp=0;

	reg state= 0;

    assign pwm_out = pwm_counter;

	always @(posedge clk) begin
        if (!resetn) begin
			counterI <= 0;
            pwm_counter <= 1;
			state<=0;
		end else begin
			counterI<= counterI+1;
            if (counterI[14] == 1) begin
				count_temp<=count_temp+1;
			end
			if (state== 1'b0 && count_temp >= pwm_in) begin
				pwm_counter<=0;
				state= 1'b1;
			end
			if (state== 1'b1 && count_temp[7] == 1) begin
				pwm_counter<=1;
				state= 1'b0;
				count_temp<=0;
			end
		end
		
	end


endmodule
